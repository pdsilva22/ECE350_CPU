module logicalA(A, B, result);
    input[31:0] A;
    input[31:0] B;
    output[31:0] result;

    and (result[0], A[0], B[0]);
    and (result[1], A[1], B[1]);
    and (result[2], A[2], B[2]);
    and (result[3], A[3], B[3]);
    and (result[4], A[4], B[4]);
    and (result[5], A[5], B[5]);
    and (result[6], A[6], B[6]);
    and (result[7], A[7], B[7]);
    and (result[8], A[8], B[8]);
    and (result[9], A[9], B[9]);
    and (result[10], A[10], B[10]);
    and (result[11], A[11], B[11]);
    and (result[12], A[12], B[12]);
    and (result[13], A[13], B[13]);
    and (result[14], A[14], B[14]);
    and (result[15], A[15], B[15]);
    and (result[16], A[16], B[16]);
    and (result[17], A[17], B[17]);
    and (result[18], A[18], B[18]);
    and (result[19], A[19], B[19]);
    and (result[20], A[20], B[20]);
    and (result[21], A[21], B[21]);
    and (result[22], A[22], B[22]);
    and (result[23], A[23], B[23]);
    and (result[24], A[24], B[24]);
    and (result[25], A[25], B[25]);
    and (result[26], A[26], B[26]);
    and (result[27], A[27], B[27]);
    and (result[28], A[28], B[28]);
    and (result[29], A[29], B[29]);
    and (result[30], A[30], B[30]);
    and (result[31], A[31], B[31]);

endmodule